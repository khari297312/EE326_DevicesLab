PreLab1
r1 2 0 100
r2 3 0 100
r3 4 0 100
r4 5 0 100
r5 6 0 100
.model BLUE D (IS = 2.659E-20 N = 2.63815 RS = 8.14349)
.model 1N4007 D  ( IS=76.9p RS=42.0m BV=1.00k IBV=5.00u
+ CJO=26.5p  M=0.333 N=1.45 TT=4.32u )
.model GREEN D (IS = 9.847E-17 N = 2.396 RS = 12.9816)
.model RED D (IS = 4.366E-25 N = 1.38167 RS = 3.00014)
.model WHITE D (IS = 1.2853E-15 N = 3.99 RS = 8.12296)
d1 1 2 1N4007
d2 1 3 BLUE
d3 1 4 GREEN
d4 1 5 RED
d5 1 6 WHITE
vin 1 0 dc 0
.dc vin 0.01 5 0.01
.control
run
plot v(2)/100 vs v(1)-v(2),v(3)/100 vs v(1)-v(3),v(4)/100 vs v(1)-v(4),v(5)/100 vs v(1)-v(5),v(6)/100 vs v(1)-v(6)
.endc
.end
