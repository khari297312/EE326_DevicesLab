RN142 PIN Diode Reverse Recovery Time
r1 2 0 100
.MODEL DRN142S D(
+ IS=127.76E-12
+ N=1.7346
+ RS=.1581
+ IKF=.14089
+ CJO=385.59E-15
+ M=.11823
+ VJ=.78827
+ ISR=139.38E-12
+ NR=3
+ BV=60
+ TT=275.00E-9)
d1 1 2 DRN142S
vin 1 0 PULSE (-1V +1V 0.02m 0.01m 0.01m 0.05m 0.1m)
.tran 0.02ms 0.2ms
.control
run
plot (v(2)/100)
plot v(1)-v(2)
.endc
.end
