Shunt Clipper DC analysis
.model d D
*r 1 3 1k
*Specifying a default diode p n
d3 0 1 d
d2 3 0 d
d1 2 1 d
d4 3 2 d

*Independent DC source whose voltage is to be varied
vin 2 0 sin (0 12v 50 0 0)

.tran 0.5ms 120ms
.control
run
*plot v(1,3)
plot v(1,3) vs v(2)
.endc
.end
