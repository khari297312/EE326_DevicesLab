.title IV Characteristics of Solar Cell

.subckt solar_cell PX NX
*IL is photo generated current (keep only 1 of the next 3 lines, whichever is necessary)
*IL NX TMP dc 0e-3    ; No light
IL NX TMP dc 10e-3   ; Illum=10mA

d1 TMP NX diode
.model diode d (is=(1e-13) n=1)

d2 TMP NX diode2
.model diode2 d (is=(2e-6) n=2)

rs TMP PX 10
rsh TMP NX 1e3

.ends solar_cell

* Define nodes
v1 N1 0 dc 0 
X1 N1 N2 solar_cell
R1 N2 0 100

* Simulation Commands
.dc v1 -2 2 0.01

.control
set TEMP=35
run
plot -i(v1) vs v(N1)-v(N2)
wrdata light_35.dat -i(v1) v(N1)-v(N2)

set TEMP=45
run
plot -i(v1) vs v(N1)-v(N2)
wrdata light_45.dat -i(v1) v(N1)-v(N2)

set TEMP=55
run
plot -i(v1) vs v(N1)-v(N2)
wrdata light_55.dat -i(v1) v(N1)-v(N2)

set TEMP=65
run
plot -i(v1) vs v(N1)-v(N2)
wrdata light_65.dat -i(v1) v(N1)-v(N2)

set TEMP=75
run
plot -i(v1) vs v(N1)-v(N2)
wrdata light_75.dat -i(v1) v(N1)-v(N2)
.endc
.end